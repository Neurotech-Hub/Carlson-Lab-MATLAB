[HEAD]:115
VPP:1.999990
OFFSET:0.000000
CHANNEL:1
RATEPOS:0.000031
RATENEG:0.000031
MAX:32767.000000
MIN:-32767.000000
[DATA]:1000
���������������������������������������������������������������������������������������������� ��������������������������������������������������������  ����������   ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������   ��������������������  ����������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������  ����������������������   ������������������������������������������������������������������������������������������������������������    ��������������  ����  
 ����������������������������������������������������������������w�\�N�I�=�&������������X�0����������L����������q�J�C�@�4�/�<�S�k��������5�d�����*�q����L�����? � � 'f��S��Q��2�%�"�d'��	�
��u��H>Nx�3�!�#=&�(�+�.I2r6;�?�BEC�?X7)j-�-�˯���{�?� ���Y�p�F�o�����������j���G � 8��C8=3,-.	
������������qXUbj`D! ( � � � � � � � � � � � � � � � � � � � � � � � { t f Z ` k i b b c \ T R R Q O Q U T F ; > H I ? 2 ) & ) , #    / 2 1 2 )      # + ,        
  ����   
 ��������  ���������������� 
   ������   ������   ��������   ���������������� ��������������������������  ���������������������������������������������������� 
 ���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� ��������������������������������������������������������������������������������������������������������������������������������������������������������  ����������������������  �������� ����������������������	  ����������������������������������  ��������